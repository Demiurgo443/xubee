module top(x0, x1, x2, x3, x4, x5, y0);
  input x0, x1, x2, x3, x4, x5;
  output y0;
  wire n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;
  assign n7 = ~x1 & ~x5;
  assign n8 = ~x2 & n7;
  assign n9 = x4 & n8;
  assign n10 = x2 & x3;
  assign n11 = n7 & ~n10;
  assign n12 = x1 & x5;
  assign n13 = x4 & ~n12;
  assign n14 = ~x3 & ~n13;
  assign n15 = x1 & x2;
  assign n16 = x5 & n15;
  assign n17 = ~x4 & n16;
  assign n18 = ~n14 & ~n17;
  assign n19 = ~n11 & n18;
  assign n20 = x0 & ~n19;
  assign n21 = x3 & ~n16;
  assign n22 = x4 & ~n15;
  assign n23 = ~n8 & ~n22;
  assign n24 = n21 & n23;
  assign n25 = ~x4 & ~x5;
  assign n26 = ~x2 ^ ~n25;
  assign n27 = ~x3 & ~n12;
  assign n28 = n26 ^ n27;
  assign n29 = x4 & x5;
  assign n30 = x2 & n29;
  assign n31 = ~n28 & ~n30;
  assign n32 = ~n24 & n31;
  assign n33 = ~x0 & ~n32;
  assign n34 = ~n20 & ~n33;
  assign n35 = ~n9 & n34;
  assign y0 = ~n35;
endmodule
