module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14;
  wire n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490;
  assign n67 = ~x0 & ~x1;
  assign n68 = x9 & ~x10;
  assign n69 = x8 & n68;
  assign n70 = x6 & n69;
  assign n71 = ~x4 & ~n70;
  assign n72 = x3 & ~n71;
  assign n73 = x2 & n72;
  assign n74 = ~x4 & ~n69;
  assign n75 = ~x3 & ~n74;
  assign n76 = x9 ^ x8;
  assign n77 = n76 ^ n68;
  assign n78 = ~x7 & ~n77;
  assign n79 = n78 ^ n68;
  assign n80 = ~x6 & n79;
  assign n81 = ~n75 & ~n80;
  assign n82 = x5 & ~n81;
  assign n83 = ~n73 & ~n82;
  assign n84 = ~n67 & ~n83;
  assign n90 = x11 & n72;
  assign n91 = x12 & ~n81;
  assign n92 = ~n90 & ~n91;
  assign n85 = ~x14 & ~n74;
  assign n86 = ~x15 & n75;
  assign n87 = ~n80 & ~n86;
  assign n88 = ~n85 & n87;
  assign n89 = x13 & ~n88;
  assign n93 = n92 ^ n89;
  assign n94 = n93 ^ n92;
  assign n95 = x16 & n72;
  assign n96 = n95 ^ n92;
  assign n97 = n96 ^ n92;
  assign n98 = ~n94 & ~n97;
  assign n99 = n98 ^ n92;
  assign n100 = n67 & n99;
  assign n101 = n100 ^ n92;
  assign n105 = x19 & ~n88;
  assign n102 = x17 & n72;
  assign n103 = x18 & ~n81;
  assign n104 = ~n102 & ~n103;
  assign n106 = n105 ^ n104;
  assign n107 = n106 ^ n104;
  assign n108 = x20 & n72;
  assign n109 = n108 ^ n104;
  assign n110 = n109 ^ n104;
  assign n111 = ~n107 & ~n110;
  assign n112 = n111 ^ n104;
  assign n113 = n67 & n112;
  assign n114 = n113 ^ n104;
  assign n118 = x23 & ~n88;
  assign n115 = x21 & n72;
  assign n116 = x22 & ~n81;
  assign n117 = ~n115 & ~n116;
  assign n119 = n118 ^ n117;
  assign n120 = n119 ^ n117;
  assign n121 = x24 & n72;
  assign n122 = n121 ^ n117;
  assign n123 = n122 ^ n117;
  assign n124 = ~n120 & ~n123;
  assign n125 = n124 ^ n117;
  assign n126 = n67 & n125;
  assign n127 = n126 ^ n117;
  assign n131 = x27 & ~n88;
  assign n128 = x25 & n72;
  assign n129 = x26 & ~n81;
  assign n130 = ~n128 & ~n129;
  assign n132 = n131 ^ n130;
  assign n133 = n132 ^ n130;
  assign n134 = x28 & n72;
  assign n135 = n134 ^ n130;
  assign n136 = n135 ^ n130;
  assign n137 = ~n133 & ~n136;
  assign n138 = n137 ^ n130;
  assign n139 = n67 & n138;
  assign n140 = n139 ^ n130;
  assign n144 = x31 & ~n88;
  assign n141 = x29 & n72;
  assign n142 = x30 & ~n81;
  assign n143 = ~n141 & ~n142;
  assign n145 = n144 ^ n143;
  assign n146 = n145 ^ n143;
  assign n147 = x32 & n72;
  assign n148 = n147 ^ n143;
  assign n149 = n148 ^ n143;
  assign n150 = ~n146 & ~n149;
  assign n151 = n150 ^ n143;
  assign n152 = n67 & n151;
  assign n153 = n152 ^ n143;
  assign n157 = x35 & ~n88;
  assign n154 = x33 & n72;
  assign n155 = x34 & ~n81;
  assign n156 = ~n154 & ~n155;
  assign n158 = n157 ^ n156;
  assign n159 = n158 ^ n156;
  assign n160 = x36 & n72;
  assign n161 = n160 ^ n156;
  assign n162 = n161 ^ n156;
  assign n163 = ~n159 & ~n162;
  assign n164 = n163 ^ n156;
  assign n165 = n67 & n164;
  assign n166 = n165 ^ n156;
  assign n167 = x37 ^ x2;
  assign n168 = ~n67 & n167;
  assign n169 = n168 ^ x2;
  assign n170 = n72 & n169;
  assign n171 = x38 ^ x5;
  assign n172 = ~n67 & n171;
  assign n173 = n172 ^ x5;
  assign n174 = ~n81 & n173;
  assign n175 = ~n170 & ~n174;
  assign n176 = ~x8 & ~x9;
  assign n177 = ~x7 & n176;
  assign n178 = x41 & ~x43;
  assign n179 = ~x42 & n178;
  assign n180 = x44 & n179;
  assign n181 = ~x42 & x43;
  assign n182 = x40 & n181;
  assign n183 = x41 & x42;
  assign n184 = ~x43 & n183;
  assign n185 = x39 & n184;
  assign n186 = ~n182 & ~n185;
  assign n187 = ~n180 & n186;
  assign n188 = n177 & ~n187;
  assign n189 = x7 & n68;
  assign n190 = ~x47 & x52;
  assign n191 = ~x46 & x48;
  assign n192 = ~n190 & ~n191;
  assign n193 = x45 & ~x51;
  assign n194 = n192 & ~n193;
  assign n195 = x49 & ~x50;
  assign n196 = ~x51 & x53;
  assign n197 = ~x52 & ~n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = x46 & ~x49;
  assign n200 = ~x45 & x50;
  assign n201 = ~n199 & ~n200;
  assign n202 = x47 & ~x48;
  assign n203 = n201 & ~n202;
  assign n204 = n198 & n203;
  assign n205 = n194 & n204;
  assign n206 = x39 & ~n205;
  assign n207 = ~x49 & ~x50;
  assign n208 = ~x51 & ~x52;
  assign n209 = x53 & n208;
  assign n210 = n207 & n209;
  assign n211 = ~x48 & n210;
  assign n212 = ~x47 & n211;
  assign n213 = ~x46 & n212;
  assign n214 = n213 ^ x45;
  assign n215 = n214 ^ n213;
  assign n216 = x50 & x51;
  assign n217 = x52 & n216;
  assign n218 = x48 & x49;
  assign n219 = n217 & n218;
  assign n220 = x47 & n219;
  assign n221 = x46 & n220;
  assign n222 = n221 ^ n213;
  assign n223 = n215 & n222;
  assign n224 = n223 ^ n213;
  assign n225 = ~x39 & n224;
  assign n226 = ~n206 & ~n225;
  assign n227 = n189 & ~n226;
  assign n228 = x8 & x9;
  assign n229 = ~x7 & n228;
  assign n230 = x44 & n229;
  assign n231 = ~n227 & ~n230;
  assign n232 = ~n188 & n231;
  assign n233 = ~x6 & ~n232;
  assign n234 = x4 & x39;
  assign n235 = n225 ^ x39;
  assign n236 = x39 ^ x7;
  assign n237 = n236 ^ x39;
  assign n238 = n235 & ~n237;
  assign n239 = n238 ^ x39;
  assign n240 = n206 ^ n70;
  assign n241 = n239 & n240;
  assign n242 = n241 ^ n206;
  assign n243 = n70 & n242;
  assign n244 = n243 ^ n70;
  assign n245 = n244 ^ n70;
  assign n246 = ~n234 & ~n245;
  assign n247 = ~n233 & n246;
  assign n248 = n247 ^ n92;
  assign n249 = ~n67 & n248;
  assign n250 = n249 ^ n92;
  assign n251 = x4 & x45;
  assign n252 = ~n67 & ~n251;
  assign n253 = ~n213 & ~n221;
  assign n254 = ~x45 & ~n253;
  assign n255 = n254 ^ x45;
  assign n256 = x45 ^ x7;
  assign n257 = n256 ^ x45;
  assign n258 = n255 & ~n257;
  assign n259 = n258 ^ x45;
  assign n260 = ~x48 & x50;
  assign n261 = n198 & ~n260;
  assign n262 = x47 & ~x49;
  assign n263 = x46 & ~x51;
  assign n264 = ~n262 & ~n263;
  assign n265 = n192 & n264;
  assign n266 = n261 & n265;
  assign n267 = x45 & ~n266;
  assign n268 = n267 ^ n70;
  assign n269 = n259 & n268;
  assign n270 = n269 ^ n267;
  assign n271 = n70 & n270;
  assign n272 = n271 ^ n70;
  assign n273 = n272 ^ n70;
  assign n274 = n252 & ~n273;
  assign n275 = n266 ^ n253;
  assign n276 = x45 & n275;
  assign n277 = n276 ^ n253;
  assign n278 = n68 & ~n277;
  assign n279 = n278 ^ x7;
  assign n280 = n279 ^ n278;
  assign n281 = x54 & n181;
  assign n282 = x45 & n184;
  assign n283 = ~n281 & ~n282;
  assign n284 = n176 & ~n283;
  assign n285 = n228 ^ x55;
  assign n286 = x10 & x56;
  assign n287 = x3 & n286;
  assign n288 = n287 ^ n228;
  assign n289 = n288 ^ n287;
  assign n290 = n176 & n179;
  assign n291 = n290 ^ n287;
  assign n292 = ~n289 & ~n291;
  assign n293 = n292 ^ n287;
  assign n294 = n285 & n293;
  assign n295 = n294 ^ x55;
  assign n296 = ~n284 & ~n295;
  assign n297 = n296 ^ n278;
  assign n298 = ~n280 & ~n297;
  assign n299 = n298 ^ n278;
  assign n300 = ~x6 & n299;
  assign n301 = n274 & ~n300;
  assign n302 = n67 & n104;
  assign n303 = ~n301 & ~n302;
  assign n305 = x51 ^ x50;
  assign n306 = x47 & ~n305;
  assign n307 = n306 ^ x50;
  assign n308 = n198 & ~n307;
  assign n309 = x52 ^ x49;
  assign n310 = ~x48 & ~n309;
  assign n311 = n310 ^ x49;
  assign n312 = n308 & n311;
  assign n304 = ~n212 & ~n220;
  assign n313 = n312 ^ n304;
  assign n314 = ~x46 & n313;
  assign n315 = n314 ^ n312;
  assign n316 = n189 & ~n315;
  assign n317 = ~n228 & ~n290;
  assign n318 = x16 & ~n317;
  assign n319 = ~x7 & n318;
  assign n320 = x13 & n181;
  assign n321 = x46 & n184;
  assign n322 = ~n320 & ~n321;
  assign n323 = n177 & ~n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = ~n316 & n324;
  assign n326 = ~x6 & ~n325;
  assign n327 = x4 & x46;
  assign n328 = ~n67 & ~n327;
  assign n329 = ~x46 & ~n304;
  assign n330 = n329 ^ x46;
  assign n331 = x46 ^ x7;
  assign n332 = n331 ^ x46;
  assign n333 = n330 & ~n332;
  assign n334 = n333 ^ x46;
  assign n335 = x46 & ~n312;
  assign n336 = n335 ^ n70;
  assign n337 = n334 & n336;
  assign n338 = n337 ^ n335;
  assign n339 = n70 & n338;
  assign n340 = n339 ^ n70;
  assign n341 = n340 ^ n70;
  assign n342 = n328 & ~n341;
  assign n343 = ~n326 & n342;
  assign n344 = n67 & n117;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~x49 & x52;
  assign n347 = x48 & ~x51;
  assign n348 = ~n346 & ~n347;
  assign n349 = n261 & n348;
  assign n350 = x47 & ~n349;
  assign n351 = ~n211 & ~n219;
  assign n352 = ~x47 & ~n351;
  assign n353 = ~n350 & ~n352;
  assign n354 = n189 & ~n353;
  assign n355 = x20 & ~n317;
  assign n356 = ~x7 & n355;
  assign n357 = x19 & n181;
  assign n358 = x47 & n184;
  assign n359 = ~n357 & ~n358;
  assign n360 = n177 & ~n359;
  assign n361 = ~n356 & ~n360;
  assign n362 = ~n354 & n361;
  assign n363 = ~x6 & ~n362;
  assign n364 = n349 ^ x47;
  assign n365 = n364 ^ n349;
  assign n366 = n351 ^ n349;
  assign n367 = ~n365 & ~n366;
  assign n368 = n367 ^ n349;
  assign n369 = ~x7 & n368;
  assign n370 = n369 ^ x47;
  assign n371 = n70 & n370;
  assign n372 = x4 & x47;
  assign n373 = ~n67 & ~n372;
  assign n374 = ~n371 & n373;
  assign n375 = ~n363 & n374;
  assign n376 = n67 & n130;
  assign n377 = ~n375 & ~n376;
  assign n378 = x49 & n217;
  assign n379 = ~x48 & n378;
  assign n380 = ~n211 & ~n379;
  assign n381 = ~n207 & ~n216;
  assign n382 = ~n197 & ~n381;
  assign n383 = ~n346 & n382;
  assign n384 = x48 & ~n383;
  assign n385 = n380 & ~n384;
  assign n386 = n189 & ~n385;
  assign n387 = x24 & ~n317;
  assign n388 = ~x7 & n387;
  assign n389 = x23 & n181;
  assign n390 = x48 & n184;
  assign n391 = ~n389 & ~n390;
  assign n392 = n177 & ~n391;
  assign n393 = ~n388 & ~n392;
  assign n394 = ~n386 & n393;
  assign n395 = ~x6 & ~n394;
  assign n396 = x4 & x48;
  assign n397 = ~n395 & ~n396;
  assign n398 = n380 ^ x48;
  assign n399 = x48 ^ x7;
  assign n400 = n399 ^ x48;
  assign n401 = ~n398 & ~n400;
  assign n402 = n401 ^ x48;
  assign n403 = n384 ^ n70;
  assign n404 = n402 & n403;
  assign n405 = n404 ^ n384;
  assign n406 = n70 & n405;
  assign n407 = n406 ^ n70;
  assign n408 = n407 ^ n70;
  assign n409 = n397 & ~n408;
  assign n410 = n409 ^ n143;
  assign n411 = ~n67 & n410;
  assign n412 = n411 ^ n143;
  assign n413 = x4 & x49;
  assign n414 = ~x50 & n208;
  assign n415 = x53 & n414;
  assign n416 = ~n217 & ~n415;
  assign n417 = x49 & n416;
  assign n418 = ~x49 & n217;
  assign n419 = ~n210 & ~n418;
  assign n420 = n419 ^ x49;
  assign n421 = ~x7 & ~n420;
  assign n422 = n421 ^ x49;
  assign n423 = ~n417 & ~n422;
  assign n424 = n70 & ~n423;
  assign n425 = ~n413 & ~n424;
  assign n426 = n425 ^ n156;
  assign n427 = n426 ^ n156;
  assign n428 = x58 & ~x63;
  assign n429 = ~x59 & ~x62;
  assign n430 = x43 & ~x61;
  assign n431 = ~x60 & n430;
  assign n432 = n429 & n431;
  assign n433 = n428 & n432;
  assign n434 = x57 & n433;
  assign n435 = n183 & n434;
  assign n436 = x27 & n181;
  assign n437 = x49 & n184;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n435 & n438;
  assign n440 = n177 & ~n439;
  assign n441 = ~n417 & n419;
  assign n442 = n189 & ~n441;
  assign n443 = x28 & ~n317;
  assign n444 = ~x7 & n443;
  assign n445 = ~n442 & ~n444;
  assign n446 = ~n440 & n445;
  assign n447 = ~x6 & ~n446;
  assign n448 = n447 ^ n156;
  assign n449 = n448 ^ n156;
  assign n450 = n427 & ~n449;
  assign n451 = n450 ^ n156;
  assign n452 = ~n67 & n451;
  assign n453 = n452 ^ n156;
  assign n457 = x32 & ~n317;
  assign n458 = ~x7 & n457;
  assign n459 = x31 & n181;
  assign n460 = x65 & n433;
  assign n461 = ~x43 & x50;
  assign n462 = x63 & x64;
  assign n463 = ~x58 & n462;
  assign n464 = n432 & n463;
  assign n465 = ~n461 & ~n464;
  assign n466 = ~n460 & n465;
  assign n467 = n183 & ~n466;
  assign n468 = ~n459 & ~n467;
  assign n469 = n177 & ~n468;
  assign n470 = ~n458 & ~n469;
  assign n471 = n196 ^ x51;
  assign n472 = ~x52 & n471;
  assign n473 = n472 ^ x51;
  assign n474 = n473 ^ x50;
  assign n475 = n189 & n474;
  assign n476 = n470 & ~n475;
  assign n477 = ~x6 & ~n476;
  assign n454 = x37 & n72;
  assign n455 = x38 & ~n81;
  assign n456 = ~n454 & ~n455;
  assign n478 = n477 ^ n456;
  assign n479 = n478 ^ n456;
  assign n480 = x4 & x50;
  assign n481 = ~x7 & n473;
  assign n482 = n481 ^ x50;
  assign n483 = n70 & n482;
  assign n484 = ~n480 & ~n483;
  assign n485 = n484 ^ n456;
  assign n486 = n485 ^ n456;
  assign n487 = ~n479 & n486;
  assign n488 = n487 ^ n456;
  assign n489 = ~n67 & n488;
  assign n490 = n489 ^ n456;
  assign y0 = n84;
  assign y1 = ~n101;
  assign y2 = ~n114;
  assign y3 = ~n127;
  assign y4 = ~n140;
  assign y5 = ~n153;
  assign y6 = ~n166;
  assign y7 = ~n175;
  assign y8 = ~n250;
  assign y9 = n303;
  assign y10 = n345;
  assign y11 = n377;
  assign y12 = ~n412;
  assign y13 = ~n453;
  assign y14 = ~n490;
endmodule
